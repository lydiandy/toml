module test

pub fn test_toml() {
}
