module toml

pub struct Encoder {
}

// the same with json.encode
pub fn encode(obj interface) ?string {
}
