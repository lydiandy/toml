module toml

pub struct Encoder {
pub mut:
	root map[string]Any
}

pub fn (mut e Encoder) encode() {
}
