module toml

//for scan each line and generate tokens
pub struct Scanner {
	text string
	pos int

}

//scan once generate one token
pub fn scan() Token {

}

pub fn (s Scanner)next() {
	
}